//------------------------------------------------------------------------
// ramtest.v
//
// This sample uses the Xilinx MIG DDR3 controller and HDL to move data
// from the PC to the DDR3 and vice-versa. Based on MIG generated example_top.v.
//
// Host Interface registers:
// WireIn 0x00
//     0 - DDR3 read enable (0=disabled, 1=enabled)
//     1 - DDR3 write enable (0=disabled, 1=enabled)
//     2 - Reset
//
// PipeIn 0x80 - DDR3 write port (U11, DDR2)
// PipeOut 0xA0 - DDR3 read port (U11, DDR2)
//
// This sample is included for reference only.  No guarantees, either
// expressed or implied, are to be drawn.
//------------------------------------------------------------------------
// tabstop 3
// Copyright (c) 2005-2016 Opal Kelly Incorporated
// $Rev$ $Date$
//------------------------------------------------------------------------
`timescale 1ns/1ps
`default_nettype none

module ramtest (
	input  wire [4:0]   okUH,
	output wire [2:0]   okHU,
	inout  wire [31:0]  okUHU,
	inout  wire         okAA,
	output wire         ok_done,

	input  wire         sys_clk_p,
	input  wire         sys_clk_n,
	
	inout  wire        si5338_scl,
	inout  wire        si5338_sda,
	
	output wire [7:0]   led,
	
	output wire         ddr4_par,     // This signal is not generated by the MIG and should be driven low
	input  wire         ddr4_alert_b, // This signal is not used by the MIG
	output wire         ddr4_ten,     // This signal is not generated by the MIG and should be driven low
	
	inout  wire [71:0]  ddr4_dq,
	inout  wire [8:0]   ddr4_dqs_t,
	inout  wire [8:0]   ddr4_dqs_c,
	inout  wire [8:0]   ddr4_dm,
	output wire [0:0]   ddr4_act_n,
	output wire [16:0]  ddr4_addr,
	output wire [1 :0]  ddr4_ba,
	output wire [0:0]   ddr4_bg,
	output wire [0 :0]  ddr4_ck_t,
	output wire [0 :0]  ddr4_ck_c,
	output wire [0 :0]  ddr4_cke,
	output wire [0 :0]  ddr4_cs_n,
	output wire [0 :0]  ddr4_odt,
	output wire         ddr4_reset_n
	);

// OK RAMTest Parameters
localparam BLOCK_SIZE = 128; // 512 bytes / 4 bytes per word, 
localparam FIFO_SIZE = 1023; // note that Xilinx does not allow use of the full 1024 words
localparam BUFFER_HEADROOM = 20; // headroom for the FIFO count to account for latency

// Capability bitfield, used to indicate features supported by this bitfile:
// [0] - Supports passing calibration status through FrontPanel
localparam CAPABILITY = 16'h0001;

wire          init_calib_complete;
reg           sys_rst;

wire [28 :0]  app_addr;
wire [2  :0]  app_cmd;
wire          app_en;
wire          app_rdy;
wire [511:0]  app_rd_data;
wire          app_rd_data_end;
wire          app_rd_data_valid;
wire [511:0]  app_wdf_data;
wire          app_wdf_end;
wire [63 :0]  app_wdf_mask;
wire          app_wdf_rdy;
wire          app_wdf_wren;

wire          clk;
wire          rst;

// Front Panel

// Target interface bus:
wire         okClk;
wire [112:0] okHE;
wire [64:0]  okEH;

wire [31:0]  ep00wire;

wire         pipe_in_read;
wire [511:0] pipe_in_data;
wire [6:0]   pipe_in_rd_count;
wire [9:0]   pipe_in_wr_count;
wire         pipe_in_valid;
wire         pipe_in_full;
wire         pipe_in_empty;
reg          pipe_in_ready;

wire         pipe_out_write;
wire [511:0] pipe_out_data;
wire [11:0]   pipe_out_rd_count;
wire [6:0]   pipe_out_wr_count;
wire         pipe_out_full;
wire         pipe_out_empty;
reg          pipe_out_ready;

// Pipe Fifos
wire         pi0_ep_write;
wire         po0_ep_read;
wire [31:0]  pi0_ep_dataout;
wire [31:0]  po0_ep_datain;

wire [63:0]  pipe_out_fifo_dout;
wire [63:0]  pipe_in_fifo_din;
reg  [ 1:0]  pipe_in_fifo_write = 2'h0;
reg  [ 1:0]  pipe_out_fifo_read = 2'h0;

assign led = {ep00wire[0],ep00wire[1],app_wdf_rdy,init_calib_complete};

	//MIG Infrastructure Reset
reg [31:0] rst_cnt;
initial rst_cnt = 32'b0;
always @(posedge okClk) begin
	if(rst_cnt < 32'h0800_0000) begin
		rst_cnt <= rst_cnt + 1;
		sys_rst <= 1'b1;
	end
	else begin
		sys_rst <= 1'b0;
	end
end

// MIG User Interface instantiation
ddr4_512_64 u_ddr4_512_64 (
  .c0_init_calib_complete(init_calib_complete),        // output wire c0_init_calib_complete
  .dbg_clk(),                                          // output wire dbg_clk
  .c0_sys_clk_p(sys_clk_p),                            // input wire c0_sys_clk_p
  .c0_sys_clk_n(sys_clk_n),                            // input wire c0_sys_clk_n
  .dbg_bus(),                                          // output wire [511 : 0] dbg_bus
  .c0_ddr4_adr(ddr4_addr),                             // output wire [16 : 0] c0_ddr4_adr
  .c0_ddr4_ba(ddr4_ba),                                // output wire [1 : 0] c0_ddr4_ba
  .c0_ddr4_cke(ddr4_cke),                              // output wire [0 : 0] c0_ddr4_cke
  .c0_ddr4_cs_n(ddr4_cs_n),                            // output wire [0 : 0] c0_ddr4_cs_n
  .c0_ddr4_dm_dbi_n(ddr4_dm),                          // inout wire [7 : 0] c0_ddr4_dm_dbi_n
  .c0_ddr4_dq(ddr4_dq),                                // inout wire [63 : 0] c0_ddr4_dq
  .c0_ddr4_dqs_c(ddr4_dqs_c),                          // inout wire [7 : 0] c0_ddr4_dqs_c
  .c0_ddr4_dqs_t(ddr4_dqs_t),                          // inout wire [7 : 0] c0_ddr4_dqs_t
  .c0_ddr4_odt(ddr4_odt),                              // output wire [0 : 0] c0_ddr4_odt
  .c0_ddr4_bg(ddr4_bg),                                // output wire [0 : 0] c0_ddr4_bg
  .c0_ddr4_reset_n(ddr4_reset_n),                      // output wire c0_ddr4_reset_n
  .c0_ddr4_act_n(ddr4_act_n),                          // output wire c0_ddr4_act_n
  .c0_ddr4_ck_c(ddr4_ck_c),                            // output wire [0 : 0] c0_ddr4_ck_c
  .c0_ddr4_ck_t(ddr4_ck_t),                            // output wire [0 : 0] c0_ddr4_ck_t

  .c0_ddr4_ui_clk(clk),               // output wire c0_ddr4_ui_clk
  .c0_ddr4_ui_clk_sync_rst(rst),      // output wire c0_ddr4_ui_clk_sync_rst
  
  .c0_ddr4_ecc_err_addr(),            // output wire [51 : 0] c0_ddr4_ecc_err_addr
  .c0_ddr4_ecc_single(),                // output wire [7 : 0] c0_ddr4_ecc_single
  .c0_ddr4_ecc_multiple(),            // output wire [7 : 0] c0_ddr4_ecc_multiple
  .c0_ddr4_app_correct_en_i(1'b1),    // input wire c0_ddr4_app_correct_en_i

  .c0_ddr4_app_en(app_en),                        // input wire c0_ddr4_app_en
  .c0_ddr4_app_hi_pri(1'b0),                // input wire c0_ddr4_app_hi_pri
  .c0_ddr4_app_wdf_end(app_wdf_end),              // input wire c0_ddr4_app_wdf_end
  .c0_ddr4_app_wdf_wren(app_wdf_wren),            // input wire c0_ddr4_app_wdf_wren
  .c0_ddr4_app_rd_data_end(app_rd_data_end),      // output wire c0_ddr4_app_rd_data_end
  .c0_ddr4_app_rd_data_valid(app_rd_data_valid),  // output wire c0_ddr4_app_rd_data_valid
  .c0_ddr4_app_rdy(app_rdy),                      // output wire c0_ddr4_app_rdy
  .c0_ddr4_app_wdf_rdy(app_wdf_rdy),              // output wire c0_ddr4_app_wdf_rdy
  .c0_ddr4_app_addr(app_addr),                    // input wire [28 : 0] c0_ddr4_app_addr
  .c0_ddr4_app_cmd(app_cmd),                      // input wire [2 : 0] c0_ddr4_app_cmd
  .c0_ddr4_app_wdf_data(app_wdf_data),            // input wire [511 : 0] c0_ddr4_app_wdf_data
  .c0_ddr4_app_wdf_mask(app_wdf_mask),            // input wire [63 : 0] c0_ddr4_app_wdf_mask
  .c0_ddr4_app_rd_data(app_rd_data),              // output wire [511 : 0] c0_ddr4_app_rd_data

  .sys_rst(sys_rst)                                      // input wire sys_rst
	);


// OK MIG DDR3 Testbench Instatiation
ddr3_test ddr3_tb (
	.clk                (clk),
	.reset              (ep00wire[2] | rst),
	.reads_en           (ep00wire[0]),
	.writes_en          (ep00wire[1]),
	.calib_done         (init_calib_complete),

	.ib_re              (pipe_in_read),
	.ib_data            (pipe_in_data),
	.ib_count           (pipe_in_rd_count),
	.ib_valid           (pipe_in_valid),
	.ib_empty           (pipe_in_empty),
	
	.ob_we              (pipe_out_write),
	.ob_data            (pipe_out_data),
	.ob_count           (pipe_out_wr_count),
	.ob_full            (pipe_out_full),
	
	.app_rdy            (app_rdy),
	.app_en             (app_en),
	.app_cmd            (app_cmd),
	.app_addr           (app_addr),
	
	.app_rd_data        (app_rd_data),
	.app_rd_data_end    (app_rd_data_end),
	.app_rd_data_valid  (app_rd_data_valid),
	
	.app_wdf_rdy        (app_wdf_rdy),
	.app_wdf_wren       (app_wdf_wren),
	.app_wdf_data       (app_wdf_data),
	.app_wdf_end        (app_wdf_end),
	.app_wdf_mask       (app_wdf_mask)
	);

//Block Throttle
always @(posedge okClk) begin
    if (sys_rst == 1'b1) begin
        pipe_in_ready <= 1'b0;
        pipe_out_ready <= 1'b0;
    end else begin
        // Check for enough space in input FIFO to pipe in another block
        // The count is compared against a reduced size to account for delays in
        // FIFO count updates.
        if(pipe_in_wr_count <= (FIFO_SIZE-BUFFER_HEADROOM-BLOCK_SIZE) ) begin
            pipe_in_ready <= 1'b1;
        end
        else begin
            pipe_in_ready <= 1'b0;
        end
    
        // Check for enough space in output FIFO to pipe out another block
        if(pipe_out_rd_count >= BLOCK_SIZE/2) begin
            pipe_out_ready <= 1'b1;
        end
        else begin
            pipe_out_ready <= 1'b0;
        end
	end
end

// Instantiate the okHost and connect endpoints.
wire [65*4-1:0]  okEHx;

okHost okHI(
	.okUH(okUH),
	.okHU(okHU),
	.okUHU(okUHU),
	.okUHs(5'b0),
	.okHUs(),
	.okUHUs(32'b0),
	.okAA(okAA),
	.okClk(okClk),
	.okHE(okHE),
	.okEH(okEH),
	.okClks(),
	.okHEs(),
	.okEHs(65'h00),
	.ok_done(ok_done)
	);

okWireOR # (.N(4)) wireOR (okEH, okEHx);
okWireIn       wi00 (.okHE(okHE),                             .ep_addr(8'h00), .ep_dataout(ep00wire));
okWireOut      wo00 (.okHE(okHE), .okEH(okEHx[ 0*65 +: 65 ]), .ep_addr(8'h20), .ep_datain({31'h00, init_calib_complete}));
okWireOut      wo01 (.okHE(okHE), .okEH(okEHx[ 1*65 +: 65 ]), .ep_addr(8'h3e), .ep_datain(CAPABILITY));
okBTPipeIn     pi0  (.okHE(okHE), .okEH(okEHx[ 2*65 +: 65 ]), .ep_addr(8'h80), .ep_write(pi0_ep_write), .ep_blockstrobe(), .ep_dataout(pi0_ep_dataout), .ep_ready(pipe_in_ready));
okBTPipeOut    po0  (.okHE(okHE), .okEH(okEHx[ 3*65 +: 65 ]), .ep_addr(8'ha0), .ep_read(po0_ep_read),   .ep_blockstrobe(), .ep_datain(po0_ep_datain),   .ep_ready(pipe_out_ready));

wire pi_translate_full, pi_translate_empty, pi_translate_valid, po_translate_full, pipe_out_valid;

fifo_w64_1024_r512_128 okPipeIn_fifo (
	.rst(ep00wire[2]),
	.wr_clk(okClk),
	.rd_clk(clk),
	.din(pipe_in_fifo_din), // Bus [63 : 0]
	.wr_en((pi_translate_valid && ~pipe_in_full)),
	.rd_en(pipe_in_read),
	.dout(pipe_in_data), // Bus [511 : 0]
	.full(pipe_in_full),
	.empty(pipe_in_empty),
	.valid(pipe_in_valid),
	.rd_data_count(pipe_in_rd_count), // Bus [6 : 0]
	.wr_data_count(pipe_in_wr_count)); // Bus [9 : 0]
	
// The Xilinx FIFO generator only translates from 512-bit down to 64-bit.
// Use a second FIFO to translate from 32-bit okPipe data to the 64-bit used
// by the Xilinx FIFO.
fifo_w32_r64 pi_translate (
  .clk(okClk),                  // input wire clk
  .srst(ep00wire[2]),                // input wire srst
  .din(pi0_ep_dataout),                  // input wire [31 : 0] din
  .wr_en(pi0_ep_write),              // input wire wr_en
  .rd_en((pi_translate_valid && ~pipe_in_full)),              // input wire rd_en
  .dout(pipe_in_fifo_din),                // output wire [63 : 0] dout
  .full(pi_translate_full),                // output wire full
  .empty(pi_translate_empty),              // output wire empty
  .valid(pi_translate_valid),
  .wr_rst_busy(),  // output wire wr_rst_busy
  .rd_rst_busy()  // output wire rd_rst_busy
);

fifo_w512_128_r64_1024 okPipeOut_fifo (
	.rst(ep00wire[2]),
	.wr_clk(clk),
	.rd_clk(okClk),
	.din(pipe_out_data), // Bus [511 : 0]
	.wr_en(pipe_out_write),
	.rd_en((~po_translate_full && pipe_out_valid)),
	.dout(pipe_out_fifo_dout), // Bus [63 : 0]
	.full(pipe_out_full),
	.empty(pipe_out_empty),
	.valid(pipe_out_valid),
	.rd_data_count(), // Bus [9 : 0]
	.wr_data_count(pipe_out_wr_count)); // Bus [6 : 0]
	
	
// The Xilinx FIFO generator only translates from 512-bit down to 64-bit.
// Use a second FIFO to translate from 32-bit okPipe data to the 64-bit used
// by the Xilinx FIFO.
fifo_w64_r32 po_translate (
  .clk(okClk),                  // input wire clk
  .srst(ep00wire[2]),                // input wire srst
  .din(pipe_out_fifo_dout),                  // input wire [31 : 0] din
  .wr_en((~po_translate_full && pipe_out_valid)),              // input wire wr_en
  .rd_en(po0_ep_read),              // input wire rd_en
  .dout(po0_ep_datain),                // output wire [63 : 0] dout
  .full(po_translate_full),                // output wire full
  .empty(),              // output wire empty
  .rd_data_count(pipe_out_rd_count)
);

endmodule
`default_nettype wire
